// connect signal to module ports

module top_module ( input a, input b, output out );
    
    mod_a instan(.in1(a),.in2(b),.out(out));

endmodule

// Create a module with one input and one output that behaves like a wire.

module top_module ( output zero );
	
	assign zero = 1'b0;
	
endmodule

// impelement out and gnd

module top_module (
    output out);
    
    assign out=1'b0;

endmodule

// impelement out and in

module top_module (
    input in,
    output out);
    assign out=in;

endmodule
